class x_sequence extends uvm_sequence;
`uvm_object_utils(x_sequence)
function new(string name = "x_sequence");
    super.new(name);
endfunction

task body;
endtask
endclass
