/* Update RTL Code Here */
/* Note : Add Commented Code and Also add summary about Code */