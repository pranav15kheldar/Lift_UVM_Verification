interface x_interface(input clk);
endinterface
