interface lift_interface(input clk);
    
endinterface
