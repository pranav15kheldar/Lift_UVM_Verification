class sequence_item extends uvm_sequence_item;
`uvm_object_utils(sequence_item)
function new(string name = "sequence_item");
    super.new(name);
endfunction

task body;
endtask
endclass
