package lift_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    `include "lift_sequence_item.sv"
    `include "lift_sequence.sv"
    `include "lift_sequencer.sv"
    `include "lift_driver.sv"
    `include "lift_monitor.sv"
    `include "lift_agent.sv"
    `include "lift_scoreboard.sv"
    `include "lift_environment.sv"
    `include "lift_test.sv"
endpackage
